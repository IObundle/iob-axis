
   ///*<InstanceName>*/
   output [7:0]  /*<InstanceName>*/_tdata,
   output        /*<InstanceName>*/_tvalid,
   input         /*<InstanceName>*/_tready,
   output        /*<InstanceName>*/_tlast,
